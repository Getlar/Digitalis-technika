`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:25:08 02/26/2019 
// Design Name: 
// Module Name:    lab2_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab2_2(
	input sw0, sw1, sw2, sw3, sw4, sw5, sw6, sw7,
	output ld0, ld1, ld2, ld3, ld4, ld5, ld6, ld7
    );
assign ld0 = sw0;
assign ld1 = sw1;
assign ld2 = sw2;
assign ld3 = sw3;
assign ld4 = sw4;
assign ld5 = sw5;
assign ld6 = sw6;
assign ld7 = sw7;


endmodule
